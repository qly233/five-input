`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   21:56:02 11/02/2021
// Design Name:   fiveinput
// Module Name:   D:/szdl/fiveinput/two.v
// Project Name:  fiveinput
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: fiveinput
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module two;

	// Inputs
	reg A;
	reg B;
	reg C;
	reg D;
	reg E;

	// Outputs
	wire F;

	// Instantiate the Unit Under Test (UUT)
	fiveinput uut (
		.A(A), 
		.B(B), 
		.C(C), 
		.D(D), 
		.E(E), 
		.F(F)
	);

	initial begin
		// Initialize Inputs
		A = 0;
		B = 0;
		C = 0;
		D = 0;
		E = 0;

		// Wait 100 ns for global reset to finish
		#100;
		A = 1;B = 0;C = 0;D = 0;E = 0;
		#100;
		A = 1;B = 1;C = 0;D = 0;E = 0;
		#100;
		A = 1;B = 1;C = 1;D = 0;E = 0;
		#100;
		A = 1;B = 0;C = 1;D = 0;E = 1;
		#100;
		A = 1;B = 0;C = 1;D = 0;E = 0;
		#100;
		A = 1;B = 0;C = 1;D = 1;E = 1;
		#100;
		A = 1;B = 1;C = 1;D = 1;E = 1;
		// Add stimulus here

	end
      
endmodule

